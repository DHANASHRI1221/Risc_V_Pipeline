// Opcode constants (subset)
`define OP_RTYPE 7'b0110011
`define OP_LOAD  7'b0000011
`define OP_STORE 7'b0100011
`define OP_BRANCH 7'b1100011