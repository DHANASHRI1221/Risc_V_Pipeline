`timescale 1ns/1ps
module write_back(input clk, input rst, input [4:0] rd_in, input [31:0] wd, input write_en);
  // This module would connect to register_file in a full design.
  // For this template, nothing is stored here.
endmodule