`timescale 1ns/1ps
// Pipeline regs placeholder: implement real fields per project needs
module pipeline_registers();
endmodule